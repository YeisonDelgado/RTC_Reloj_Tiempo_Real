-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Wed Dec 14 21:33:43 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Display7seg IS 
	PORT
	(
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		C1 :  IN  STD_LOGIC;
		D1 :  IN  STD_LOGIC;
		a :  OUT  STD_LOGIC;
		b :  OUT  STD_LOGIC;
		c :  OUT  STD_LOGIC;
		d :  OUT  STD_LOGIC;
		e :  OUT  STD_LOGIC;
		f :  OUT  STD_LOGIC;
		g :  OUT  STD_LOGIC
	);
END Display7seg;

ARCHITECTURE bdf_type OF Display7seg IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_47 <= NOT(D1 XOR B1);


SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_0 AND C1;


SYNTHESIZED_WIRE_1 <= NOT(C1 XOR D1);


SYNTHESIZED_WIRE_39 <= A1 OR SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_46;


SYNTHESIZED_WIRE_35 <= A1 OR SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_51 <= NOT(C1);



SYNTHESIZED_WIRE_11 <= NOT(A1);



SYNTHESIZED_WIRE_38 <= A1 OR SYNTHESIZED_WIRE_47 OR C1;


SYNTHESIZED_WIRE_12 <= NOT(B1);



SYNTHESIZED_WIRE_48 <= NOT(C1);



SYNTHESIZED_WIRE_29 <= NOT(A1);



SYNTHESIZED_WIRE_50 <= NOT(B1);



SYNTHESIZED_WIRE_49 <= NOT(D1);



SYNTHESIZED_WIRE_40 <= A1 OR SYNTHESIZED_WIRE_48 OR D1 OR B1;


SYNTHESIZED_WIRE_42 <= SYNTHESIZED_WIRE_49 AND SYNTHESIZED_WIRE_8;


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_46 <= SYNTHESIZED_WIRE_11 AND SYNTHESIZED_WIRE_12;


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_50 AND SYNTHESIZED_WIRE_51;


SYNTHESIZED_WIRE_44 <= SYNTHESIZED_WIRE_51 OR SYNTHESIZED_WIRE_16;


SYNTHESIZED_WIRE_34 <= A1 OR SYNTHESIZED_WIRE_17 OR SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_23 <= NOT(D1);



SYNTHESIZED_WIRE_43 <= NOT(C1);



SYNTHESIZED_WIRE_45 <= SYNTHESIZED_WIRE_46 OR SYNTHESIZED_WIRE_20;


SYNTHESIZED_WIRE_20 <= NOT(D1);



SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_16 <= C1 AND SYNTHESIZED_WIRE_23;


SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_24 AND SYNTHESIZED_WIRE_48;


SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27;


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_28 AND A1;


SYNTHESIZED_WIRE_28 <= NOT(D1);



SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_29 AND SYNTHESIZED_WIRE_50;


SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_33 AND C1;


SYNTHESIZED_WIRE_0 <= NOT(A1);



f <= NOT(SYNTHESIZED_WIRE_34);



g <= NOT(SYNTHESIZED_WIRE_35);



SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_49 AND SYNTHESIZED_WIRE_51;


a <= NOT(SYNTHESIZED_WIRE_38);



b <= NOT(SYNTHESIZED_WIRE_39);



c <= NOT(SYNTHESIZED_WIRE_40);



d <= NOT(SYNTHESIZED_WIRE_41);



e <= NOT(SYNTHESIZED_WIRE_42);



SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_43 AND B1;


SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_44 AND B1;


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_45 AND C1;


END bdf_type;